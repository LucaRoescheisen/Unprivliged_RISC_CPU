module top();




endmodule